module SFRReader(  
    input clk,
    input [7:0] addr,
    output [7:0] val,
);

endmodule