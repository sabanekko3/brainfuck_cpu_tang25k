module SFRWriter(  
    input clk,
    input [7:0] val,
    input [7:0] addr,
    input valid
);

endmodule