module ROM (
    input [7:0] addr,
    output reg [2:0] code,
    output rom_overrun
);
`define INC  3'b111 //+
`define DEC  3'b110 //-
`define MOVR 3'b101 //>
`define MOVL 3'b100 //<
`define IF   3'b011 //[
`define BACK 3'b010 //]
`define OUT  3'b001 //.
`define NOP  3'b000 //,

localparam len = 124;

 wire [2:0] rom_array[0:len-1] = '{
    `DEC,
    `DEC,
    `IF,
    `DEC,
    `DEC,
    `DEC,
    `DEC,
    `DEC,
    `MOVR,
    `INC,
    `MOVL,
    `BACK,
    `MOVR,
    `DEC,
    `DEC,
    `DEC,
    `DEC,
    `OUT,
    `IF,
    `DEC,
    `DEC,
    `DEC,
    `MOVR,
    `INC,
    `MOVL,
    `BACK,
    `MOVR,
    `DEC,
    `DEC,
    `DEC,
    `DEC,
    `OUT,
    `INC,
    `INC,
    `INC,
    `IF,
    `DEC,
    `MOVR,
    `INC,
    `INC,
    `INC,
    `MOVL,
    `BACK,
    `MOVR,
    `INC,
    `INC,
    `OUT,
    `INC,
    `INC,
    `INC,
    `INC,
    `INC,
    `INC,
    `INC,
    `INC,
    `OUT,
    `INC,
    `INC,
    `INC,
    `INC,
    `INC,
    `OUT,
    `DEC,
    `IF,
    `DEC,
    `MOVR,
    `INC,
    `INC,
    `INC,
    `MOVL,
    `BACK,
    `MOVR,
    `DEC,
    `OUT,
    `MOVR,
    `DEC,
    `IF,
    `DEC,
    `DEC,
    `DEC,
    `MOVR,
    `INC,
    `MOVL,
    `BACK,
    `MOVR,
    `OUT,
    `DEC,
    `IF,
    `DEC,
    `DEC,
    `DEC,
    `DEC,
    `DEC,
    `MOVR,
    `INC,
    `MOVL,
    `BACK,
    `MOVR,
    `DEC,
    `OUT,
    `INC,
    `INC,
    `INC,
    `INC,
    `INC,
    `INC,
    `INC,
    `INC,
    `OUT,
    `DEC,
    `IF,
    `DEC,
    `DEC,
    `MOVR,
    `INC,
    `MOVL,
    `BACK,
    `MOVR,
    `DEC,
    `DEC,
    `DEC,
    `DEC,
    `OUT,
    `OUT
};

assign code = addr < len ? rom_array[addr] : 3'h0;
assign rom_overrun =  addr < len ? 1'h0 : 1'h1;

endmodule
