module ROM (
    input [9:0] addr,
    output reg [2:0] code,
    output rom_overrun
);
`define INC  3'b111 //+
`define DEC  3'b110 //-
`define MOVR 3'b101 //>
`define MOVL 3'b100 //<
`define IF   3'b011 //[
`define BACK 3'b010 //]
`define OUT  3'b001 //.
`define IN  3'b000 //,

localparam len = 470;

always_comb begin
    case(addr)
        10'h000:code <= `MOVR;
        10'h001:code <= `MOVR;
        10'h002:code <= `INC;
        10'h003:code <= `MOVR;
        10'h004:code <= `INC;
        10'h005:code <= `INC;
        10'h006:code <= `INC;
        10'h007:code <= `INC;
        10'h008:code <= `INC;
        10'h009:code <= `INC;
        10'h00a:code <= `INC;
        10'h00b:code <= `INC;
        10'h00c:code <= `INC;
        10'h00d:code <= `INC;
        10'h00e:code <= `INC;
        10'h00f:code <= `INC;
        10'h010:code <= `OUT;
        10'h011:code <= `MOVR;
        10'h012:code <= `MOVR;
        10'h013:code <= `INC;
        10'h014:code <= `INC;
        10'h015:code <= `INC;
        10'h016:code <= `INC;
        10'h017:code <= `INC;
        10'h018:code <= `INC;
        10'h019:code <= `INC;
        10'h01a:code <= `INC;
        10'h01b:code <= `MOVR;
        10'h01c:code <= `INC;
        10'h01d:code <= `INC;
        10'h01e:code <= `INC;
        10'h01f:code <= `INC;
        10'h020:code <= `INC;
        10'h021:code <= `INC;
        10'h022:code <= `INC;
        10'h023:code <= `INC;
        10'h024:code <= `MOVR;
        10'h025:code <= `INC;
        10'h026:code <= `MOVR;
        10'h027:code <= `MOVR;
        10'h028:code <= `MOVR;
        10'h029:code <= `INC;
        10'h02a:code <= `MOVR;
        10'h02b:code <= `MOVR;
        10'h02c:code <= `MOVR;
        10'h02d:code <= `MOVL;
        10'h02e:code <= `MOVL;
        10'h02f:code <= `MOVL;
        10'h030:code <= `MOVL;
        10'h031:code <= `MOVL;
        10'h032:code <= `MOVL;
        10'h033:code <= `MOVL;
        10'h034:code <= `MOVL;
        10'h035:code <= `MOVL;
        10'h036:code <= `MOVL;
        10'h037:code <= `MOVL;
        10'h038:code <= `IF;
        10'h039:code <= `MOVR;
        10'h03a:code <= `MOVR;
        10'h03b:code <= `MOVR;
        10'h03c:code <= `MOVR;
        10'h03d:code <= `MOVR;
        10'h03e:code <= `MOVR;
        10'h03f:code <= `INC;
        10'h040:code <= `MOVL;
        10'h041:code <= `IF;
        10'h042:code <= `MOVL;
        10'h043:code <= `MOVL;
        10'h044:code <= `MOVL;
        10'h045:code <= `INC;
        10'h046:code <= `OUT;
        10'h047:code <= `MOVR;
        10'h048:code <= `MOVR;
        10'h049:code <= `MOVR;
        10'h04a:code <= `MOVR;
        10'h04b:code <= `DEC;
        10'h04c:code <= `BACK;
        10'h04d:code <= `MOVR;
        10'h04e:code <= `IF;
        10'h04f:code <= `DEC;
        10'h050:code <= `MOVL;
        10'h051:code <= `MOVL;
        10'h052:code <= `MOVL;
        10'h053:code <= `MOVL;
        10'h054:code <= `DEC;
        10'h055:code <= `OUT;
        10'h056:code <= `MOVR;
        10'h057:code <= `MOVR;
        10'h058:code <= `MOVR;
        10'h059:code <= `MOVR;
        10'h05a:code <= `MOVR;
        10'h05b:code <= `BACK;
        10'h05c:code <= `MOVL;
        10'h05d:code <= `INC;
        10'h05e:code <= `MOVL;
        10'h05f:code <= `MOVL;
        10'h060:code <= `MOVL;
        10'h061:code <= `MOVL;
        10'h062:code <= `IF;
        10'h063:code <= `MOVR;
        10'h064:code <= `MOVR;
        10'h065:code <= `MOVR;
        10'h066:code <= `MOVR;
        10'h067:code <= `DEC;
        10'h068:code <= `BACK;
        10'h069:code <= `MOVR;
        10'h06a:code <= `MOVR;
        10'h06b:code <= `MOVR;
        10'h06c:code <= `MOVR;
        10'h06d:code <= `IF;
        10'h06e:code <= `DEC;
        10'h06f:code <= `MOVL;
        10'h070:code <= `INC;
        10'h071:code <= `MOVR;
        10'h072:code <= `MOVR;
        10'h073:code <= `MOVR;
        10'h074:code <= `MOVR;
        10'h075:code <= `MOVR;
        10'h076:code <= `BACK;
        10'h077:code <= `MOVL;
        10'h078:code <= `MOVL;
        10'h079:code <= `MOVL;
        10'h07a:code <= `MOVL;
        10'h07b:code <= `INC;
        10'h07c:code <= `MOVL;
        10'h07d:code <= `MOVL;
        10'h07e:code <= `MOVL;
        10'h07f:code <= `MOVL;
        10'h080:code <= `DEC;
        10'h081:code <= `DEC;
        10'h082:code <= `DEC;
        10'h083:code <= `DEC;
        10'h084:code <= `DEC;
        10'h085:code <= `DEC;
        10'h086:code <= `DEC;
        10'h087:code <= `DEC;
        10'h088:code <= `DEC;
        10'h089:code <= `DEC;
        10'h08a:code <= `DEC;
        10'h08b:code <= `DEC;
        10'h08c:code <= `IF;
        10'h08d:code <= `MOVR;
        10'h08e:code <= `MOVR;
        10'h08f:code <= `MOVR;
        10'h090:code <= `MOVR;
        10'h091:code <= `DEC;
        10'h092:code <= `BACK;
        10'h093:code <= `MOVR;
        10'h094:code <= `MOVR;
        10'h095:code <= `MOVR;
        10'h096:code <= `MOVR;
        10'h097:code <= `IF;
        10'h098:code <= `DEC;
        10'h099:code <= `MOVL;
        10'h09a:code <= `DEC;
        10'h09b:code <= `MOVR;
        10'h09c:code <= `MOVR;
        10'h09d:code <= `MOVR;
        10'h09e:code <= `MOVR;
        10'h09f:code <= `MOVR;
        10'h0a0:code <= `BACK;
        10'h0a1:code <= `MOVL;
        10'h0a2:code <= `MOVL;
        10'h0a3:code <= `MOVL;
        10'h0a4:code <= `MOVL;
        10'h0a5:code <= `MOVL;
        10'h0a6:code <= `MOVL;
        10'h0a7:code <= `MOVL;
        10'h0a8:code <= `MOVL;
        10'h0a9:code <= `INC;
        10'h0aa:code <= `INC;
        10'h0ab:code <= `INC;
        10'h0ac:code <= `INC;
        10'h0ad:code <= `INC;
        10'h0ae:code <= `INC;
        10'h0af:code <= `INC;
        10'h0b0:code <= `INC;
        10'h0b1:code <= `INC;
        10'h0b2:code <= `INC;
        10'h0b3:code <= `INC;
        10'h0b4:code <= `INC;
        10'h0b5:code <= `MOVL;
        10'h0b6:code <= `MOVL;
        10'h0b7:code <= `MOVR;
        10'h0b8:code <= `MOVR;
        10'h0b9:code <= `MOVR;
        10'h0ba:code <= `MOVR;
        10'h0bb:code <= `MOVR;
        10'h0bc:code <= `MOVR;
        10'h0bd:code <= `MOVR;
        10'h0be:code <= `MOVR;
        10'h0bf:code <= `MOVR;
        10'h0c0:code <= `INC;
        10'h0c1:code <= `MOVL;
        10'h0c2:code <= `IF;
        10'h0c3:code <= `MOVL;
        10'h0c4:code <= `MOVL;
        10'h0c5:code <= `MOVL;
        10'h0c6:code <= `MOVL;
        10'h0c7:code <= `MOVL;
        10'h0c8:code <= `INC;
        10'h0c9:code <= `OUT;
        10'h0ca:code <= `MOVR;
        10'h0cb:code <= `MOVR;
        10'h0cc:code <= `MOVR;
        10'h0cd:code <= `MOVR;
        10'h0ce:code <= `MOVR;
        10'h0cf:code <= `MOVR;
        10'h0d0:code <= `DEC;
        10'h0d1:code <= `BACK;
        10'h0d2:code <= `MOVR;
        10'h0d3:code <= `IF;
        10'h0d4:code <= `DEC;
        10'h0d5:code <= `MOVL;
        10'h0d6:code <= `MOVL;
        10'h0d7:code <= `MOVL;
        10'h0d8:code <= `MOVL;
        10'h0d9:code <= `MOVL;
        10'h0da:code <= `MOVL;
        10'h0db:code <= `DEC;
        10'h0dc:code <= `OUT;
        10'h0dd:code <= `MOVR;
        10'h0de:code <= `MOVR;
        10'h0df:code <= `MOVR;
        10'h0e0:code <= `MOVR;
        10'h0e1:code <= `MOVR;
        10'h0e2:code <= `MOVR;
        10'h0e3:code <= `MOVR;
        10'h0e4:code <= `BACK;
        10'h0e5:code <= `MOVL;
        10'h0e6:code <= `MOVL;
        10'h0e7:code <= `MOVL;
        10'h0e8:code <= `MOVL;
        10'h0e9:code <= `INC;
        10'h0ea:code <= `MOVL;
        10'h0eb:code <= `MOVL;
        10'h0ec:code <= `MOVL;
        10'h0ed:code <= `IF;
        10'h0ee:code <= `MOVR;
        10'h0ef:code <= `MOVR;
        10'h0f0:code <= `MOVR;
        10'h0f1:code <= `DEC;
        10'h0f2:code <= `BACK;
        10'h0f3:code <= `MOVR;
        10'h0f4:code <= `MOVR;
        10'h0f5:code <= `MOVR;
        10'h0f6:code <= `IF;
        10'h0f7:code <= `DEC;
        10'h0f8:code <= `MOVR;
        10'h0f9:code <= `MOVR;
        10'h0fa:code <= `INC;
        10'h0fb:code <= `MOVR;
        10'h0fc:code <= `BACK;
        10'h0fd:code <= `MOVL;
        10'h0fe:code <= `MOVL;
        10'h0ff:code <= `MOVL;
        10'h100:code <= `INC;
        10'h101:code <= `MOVL;
        10'h102:code <= `MOVL;
        10'h103:code <= `MOVL;
        10'h104:code <= `DEC;
        10'h105:code <= `DEC;
        10'h106:code <= `DEC;
        10'h107:code <= `DEC;
        10'h108:code <= `DEC;
        10'h109:code <= `DEC;
        10'h10a:code <= `DEC;
        10'h10b:code <= `DEC;
        10'h10c:code <= `DEC;
        10'h10d:code <= `DEC;
        10'h10e:code <= `DEC;
        10'h10f:code <= `DEC;
        10'h110:code <= `IF;
        10'h111:code <= `MOVR;
        10'h112:code <= `MOVR;
        10'h113:code <= `MOVR;
        10'h114:code <= `DEC;
        10'h115:code <= `BACK;
        10'h116:code <= `MOVR;
        10'h117:code <= `MOVR;
        10'h118:code <= `MOVR;
        10'h119:code <= `IF;
        10'h11a:code <= `DEC;
        10'h11b:code <= `MOVR;
        10'h11c:code <= `MOVR;
        10'h11d:code <= `DEC;
        10'h11e:code <= `MOVR;
        10'h11f:code <= `BACK;
        10'h120:code <= `MOVL;
        10'h121:code <= `MOVL;
        10'h122:code <= `MOVL;
        10'h123:code <= `MOVL;
        10'h124:code <= `MOVL;
        10'h125:code <= `MOVL;
        10'h126:code <= `INC;
        10'h127:code <= `INC;
        10'h128:code <= `INC;
        10'h129:code <= `INC;
        10'h12a:code <= `INC;
        10'h12b:code <= `INC;
        10'h12c:code <= `INC;
        10'h12d:code <= `INC;
        10'h12e:code <= `INC;
        10'h12f:code <= `INC;
        10'h130:code <= `INC;
        10'h131:code <= `INC;
        10'h132:code <= `MOVL;
        10'h133:code <= `MOVL;
        10'h134:code <= `MOVL;
        10'h135:code <= `MOVR;
        10'h136:code <= `MOVR;
        10'h137:code <= `MOVR;
        10'h138:code <= `MOVR;
        10'h139:code <= `MOVR;
        10'h13a:code <= `MOVR;
        10'h13b:code <= `MOVR;
        10'h13c:code <= `MOVR;
        10'h13d:code <= `MOVR;
        10'h13e:code <= `MOVR;
        10'h13f:code <= `MOVR;
        10'h140:code <= `MOVR;
        10'h141:code <= `INC;
        10'h142:code <= `MOVL;
        10'h143:code <= `IF;
        10'h144:code <= `MOVL;
        10'h145:code <= `MOVL;
        10'h146:code <= `MOVL;
        10'h147:code <= `MOVL;
        10'h148:code <= `MOVL;
        10'h149:code <= `MOVL;
        10'h14a:code <= `MOVL;
        10'h14b:code <= `INC;
        10'h14c:code <= `OUT;
        10'h14d:code <= `MOVR;
        10'h14e:code <= `MOVR;
        10'h14f:code <= `MOVR;
        10'h150:code <= `MOVR;
        10'h151:code <= `MOVR;
        10'h152:code <= `MOVR;
        10'h153:code <= `MOVR;
        10'h154:code <= `MOVR;
        10'h155:code <= `DEC;
        10'h156:code <= `BACK;
        10'h157:code <= `MOVR;
        10'h158:code <= `IF;
        10'h159:code <= `DEC;
        10'h15a:code <= `MOVL;
        10'h15b:code <= `MOVL;
        10'h15c:code <= `MOVL;
        10'h15d:code <= `MOVL;
        10'h15e:code <= `MOVL;
        10'h15f:code <= `MOVL;
        10'h160:code <= `MOVL;
        10'h161:code <= `MOVL;
        10'h162:code <= `DEC;
        10'h163:code <= `OUT;
        10'h164:code <= `MOVR;
        10'h165:code <= `MOVR;
        10'h166:code <= `MOVR;
        10'h167:code <= `MOVR;
        10'h168:code <= `MOVR;
        10'h169:code <= `MOVR;
        10'h16a:code <= `MOVR;
        10'h16b:code <= `MOVR;
        10'h16c:code <= `MOVR;
        10'h16d:code <= `BACK;
        10'h16e:code <= `MOVL;
        10'h16f:code <= `MOVL;
        10'h170:code <= `MOVL;
        10'h171:code <= `MOVL;
        10'h172:code <= `INC;
        10'h173:code <= `MOVL;
        10'h174:code <= `MOVL;
        10'h175:code <= `MOVL;
        10'h176:code <= `MOVL;
        10'h177:code <= `MOVL;
        10'h178:code <= `IF;
        10'h179:code <= `MOVR;
        10'h17a:code <= `MOVR;
        10'h17b:code <= `MOVR;
        10'h17c:code <= `MOVR;
        10'h17d:code <= `MOVR;
        10'h17e:code <= `DEC;
        10'h17f:code <= `BACK;
        10'h180:code <= `MOVR;
        10'h181:code <= `MOVR;
        10'h182:code <= `MOVR;
        10'h183:code <= `MOVR;
        10'h184:code <= `MOVR;
        10'h185:code <= `IF;
        10'h186:code <= `DEC;
        10'h187:code <= `MOVR;
        10'h188:code <= `MOVR;
        10'h189:code <= `INC;
        10'h18a:code <= `MOVR;
        10'h18b:code <= `MOVR;
        10'h18c:code <= `MOVR;
        10'h18d:code <= `BACK;
        10'h18e:code <= `MOVL;
        10'h18f:code <= `MOVL;
        10'h190:code <= `MOVL;
        10'h191:code <= `MOVL;
        10'h192:code <= `MOVL;
        10'h193:code <= `INC;
        10'h194:code <= `MOVL;
        10'h195:code <= `MOVL;
        10'h196:code <= `MOVL;
        10'h197:code <= `MOVL;
        10'h198:code <= `MOVL;
        10'h199:code <= `DEC;
        10'h19a:code <= `DEC;
        10'h19b:code <= `DEC;
        10'h19c:code <= `DEC;
        10'h19d:code <= `DEC;
        10'h19e:code <= `DEC;
        10'h19f:code <= `DEC;
        10'h1a0:code <= `DEC;
        10'h1a1:code <= `DEC;
        10'h1a2:code <= `DEC;
        10'h1a3:code <= `DEC;
        10'h1a4:code <= `DEC;
        10'h1a5:code <= `IF;
        10'h1a6:code <= `MOVR;
        10'h1a7:code <= `MOVR;
        10'h1a8:code <= `MOVR;
        10'h1a9:code <= `MOVR;
        10'h1aa:code <= `MOVR;
        10'h1ab:code <= `DEC;
        10'h1ac:code <= `BACK;
        10'h1ad:code <= `MOVR;
        10'h1ae:code <= `MOVR;
        10'h1af:code <= `MOVR;
        10'h1b0:code <= `MOVR;
        10'h1b1:code <= `MOVR;
        10'h1b2:code <= `IF;
        10'h1b3:code <= `DEC;
        10'h1b4:code <= `MOVR;
        10'h1b5:code <= `MOVR;
        10'h1b6:code <= `DEC;
        10'h1b7:code <= `MOVR;
        10'h1b8:code <= `MOVR;
        10'h1b9:code <= `MOVR;
        10'h1ba:code <= `BACK;
        10'h1bb:code <= `MOVL;
        10'h1bc:code <= `MOVL;
        10'h1bd:code <= `MOVL;
        10'h1be:code <= `MOVL;
        10'h1bf:code <= `MOVL;
        10'h1c0:code <= `MOVL;
        10'h1c1:code <= `MOVL;
        10'h1c2:code <= `MOVL;
        10'h1c3:code <= `MOVL;
        10'h1c4:code <= `MOVL;
        10'h1c5:code <= `INC;
        10'h1c6:code <= `INC;
        10'h1c7:code <= `INC;
        10'h1c8:code <= `INC;
        10'h1c9:code <= `INC;
        10'h1ca:code <= `INC;
        10'h1cb:code <= `INC;
        10'h1cc:code <= `INC;
        10'h1cd:code <= `INC;
        10'h1ce:code <= `INC;
        10'h1cf:code <= `INC;
        10'h1d0:code <= `INC;
        10'h1d1:code <= `MOVL;
        10'h1d2:code <= `MOVL;
        10'h1d3:code <= `MOVL;
        10'h1d4:code <= `MOVL;
        10'h1d5:code <= `BACK;
        default:code <=  `INC;
    endcase
end

assign rom_overrun =  addr < len ? 1'h0 : 1'h1;

endmodule
